/*
 Message Types
 Author: Hyoukjun Kwon(hyoukjun@gatech.edu)

*/


/********** Native Libraries ************/
import Vector::*;
/******** User-Defined Libraries *********/
import NetworkTypes::*;
import VirtualChannelTypes::*;
import RoutingTypes::*;

/************* Definitions **************/

//1. Sub-definitions for Flit class
  //Message class and Flit types
  typedef Data FlitData;

  // Flit Type
  typedef struct {
    FlitType flitType;    // Identify the type of flit: Head, Body, Tail
    FlitData  flitData;   // The actual data.
  } Flit deriving (Bits, Eq);

  instance FShow#(Flit);
    function Fmt fshow (Flit flit);
        return ($format("<Flit:")
                +
                $format("\tFlitType(%0d)>", flit.flitType)
                +
                $format("\tFlitData(%0h)", flit.flitData)
                );
    endfunction
  endinstance

  typedef struct {
    Flit flit;        // Actual Router Flit
    DirIdx destDirn;  // Output port in current switch: To be generated by Route Computation Unit
  } SwitchFlit deriving (Bits, Eq);

  instance FShow#(SwitchFlit);
    function Fmt fshow (SwitchFlit switchFlit);
        return ($format("<SwitchFlit:")
                +
                $format("SwitchDirection(%0d)", switchFlit.destDirn)
                +
                $format("\tFlit(%s)>", fshow(switchFlit.flit))
                );
    endfunction
  endinstance

/* Bundles */
// typedef Vector#(NumPorts, Maybe#(Header))   HeaderBundle;
typedef Vector#(NumPorts, Flit)     FlitBundle;

