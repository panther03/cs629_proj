import Core::*;
module mkTopPipelined(Empty);
    Core core <- mkCore(0);
endmodule
